`default_nettype none

module moduleName (
    ports
);


endmodule